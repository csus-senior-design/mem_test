
module ISSP (
	probe,
	source_clk,
	source);	

	input	[1:0]	probe;
	input		source_clk;
	output	[2:0]	source;
endmodule
